module STOPWATCH_tb;

reg CLK;
wire [3:0] HOUR;
wire [2:0] MINHIGH;
wire [3:0] MINLOW;
wire [3:0] MSE00;
wire [3:0] MSEC1ST;
wire [3:0] MSEC2ND;
reg RST;
wire [2:0] SECHIGH;
wire [3:0] SECLOW;
reg STOPWATCH_RUN;
reg SW_F1;
reg SW_F2;

STOPWATCH
 U0 (
  .CLK(CLK),
  .HOUR(HOUR),
  .MINHIGH(MINHIGH),
  .MINLOW(MINLOW),
  .MSE00(MSE00),
  .MSEC1ST(MSEC1ST),
  .MSEC2ND(MSEC2ND),
  .RST(RST),
  .SECHIGH(SECHIGH),
  .SECLOW(SECLOW),
  .STOPWATCH_RUN(STOPWATCH_RUN),
  .SW_F1(SW_F1),
  .SW_F2(SW_F2));

  initial
  begin
    CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
    #100 CLK = 1'b0;
    #100 CLK = 1'b1;
  end

  initial
  begin
    RST = 1'b0;
    #100 RST = 1'b1;
    #200 RST = 1'b0;
  end

  initial
  begin
    STOPWATCH_RUN = 1'b0;
    #400 STOPWATCH_RUN = 1'b1;
  end

  initial
  begin
    SW_F1 = 1'b0;
    #600 SW_F1 = 1'b1;
    #300 SW_F1 = 1'b0;
    #2200 SW_F1 = 1'b1;
    #200 SW_F1 = 1'b0;
  end

  initial
  begin
    SW_F2 = 1'b0;
    #3700 SW_F2 = 1'b1;
    #200 SW_F2 = 1'b0;
  end

endmodule
