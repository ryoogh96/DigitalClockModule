module conticonti(p00,p01,p02,p03,p04,p05,p06,p07,p08,p09,p10,p11,p12,p13,p14,p15,p16,p17,p18,p19,p20,p21,p22,p23,p24,p25,p26,p27,p28,p29,p30,p31,p32,p33,p34,p35,p36,p37,p38,p39,p40,p41,p42,p43,p44,p45,p46,p47,p48,p49,p50,p51,p52,p53,p54,p55,p56,p57,p58,p59,p60,p61,p62,p63);

input p00;
input p01;
input p02;
input p03;
input p04;
input p05;
input p06;
input p07;
input p08;
input p09;
input p10;
input p11;
input p12;
input p13;
input p14;
input p15;
input p16;
input p17;
input p18;
input p19;
input p20;
input p21;
input p22;
input p23;
input p24;
input p25;
input p26;
input p27;
input p28;
input p29;
input p30;
input p31;
output p32;
output p33;
output p34;
output p35;
output p36;
output p37;
output p38;
output p39;
output p40;
output p41;
output p42;
output p43;
output p44;
output p45;
output p46;
output p47;
output p48;
output p49;
output p50;
output p51;
output p52;
output p53;
output p54;
output p55;
output p56;
output p57;
output p58;
output p59;
output p60;
output p61;
output p62;
output p63;

wire  w0;
wire  w1;
wire  w2;
wire  w3;
wire  w4;
wire  w5;
wire  w6;
wire  w7;
wire  w8;
wire  w9;
wire  w10;
wire  w11;
wire  w12;
wire  w13;
wire  w14;
wire  w15;
wire  w16;
wire  w17;
wire  w18;
wire  w19;
wire  w20;
wire  w21;
wire  w22;
wire  w23;
wire  w24;
wire  w25;
wire  w26;
wire  w27;
wire  w28;
wire  w29;
wire  w30;
wire  w31;

assign w0 = p00;
assign w1 = p01;
assign w2 = p02;
assign w3 = p03;
assign w4 = p04;
assign w5 = p05;
assign w6 = p06;
assign w7 = p07;
assign w8 = p08;
assign w9 = p09;
assign w10 = p10;
assign w11 = p11;
assign w12 = p12;
assign w13 = p13;
assign w14 = p14;
assign w15 = p15;
assign w16 = p16;
assign w17 = p17;
assign w18 = p18;
assign w19 = p19;
assign w20 = p20;
assign w21 = p21;
assign w22 = p22;
assign w23 = p23;
assign w24 = p24;
assign w25 = p25;
assign w26 = p26;
assign w27 = p27;
assign w28 = p28;
assign w29 = p29;
assign w30 = p30;
assign w31 = p31;
assign p32 = w0;
assign p33 = w1;
assign p34 = w2;
assign p35 = w3;
assign p36 = w4;
assign p37 = w5;
assign p38 = w6;
assign p39 = w7;
assign p40 = w8;
assign p41 = w9;
assign p42 = w10;
assign p43 = w11;
assign p44 = w12;
assign p45 = w13;
assign p46 = w14;
assign p47 = w15;
assign p48 = w16;
assign p49 = w17;
assign p50 = w18;
assign p51 = w19;
assign p52 = w20;
assign p53 = w21;
assign p54 = w22;
assign p55 = w23;
assign p56 = w24;
assign p57 = w25;
assign p58 = w26;
assign p59 = w27;
assign p60 = w28;
assign p61 = w29;
assign p62 = w30;
assign p63 = w31;

endmodule

