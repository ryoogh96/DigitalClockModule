module counter60to7seg_tb;

wire [6:0] HOUR1;
wire [6:0] HOUR10;
wire [6:0] MIN1;
wire [6:0] MIN10;
wire [6:0] SEC1;
wire [6:0] SEC10;
reg clk;
reg rst;

counter60to7seg
 U0 (
  .HOUR1(HOUR1),
  .HOUR10(HOUR10),
  .MIN1(MIN1),
  .MIN10(MIN10),
  .SEC1(SEC1),
  .SEC10(SEC10),
  .clk(clk),
  .rst(rst));

  initial
  begin
    clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
    #10 clk = 1'b1;
    #10 clk = 1'b0;
  end

  initial
  begin
    rst = 1'b0;
    #100 rst = 1'b1;
    #100 rst = 1'b0;
  end

endmodule
